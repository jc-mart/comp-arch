`define arithmetic_base 32'bxxxxxxxxxxxxxxxxxxxxxxxxx0110011
`define arithmetic_imm  32'bxxxxxxxxxxxxxxxxxxxxxxxxx0010011
`define load            32'bxxxxxxxxxxxxxxxxxxxxxxxxx0000011
`define store           32'bxxxxxxxxxxxxxxxxxxxxxxxxx0100011
`define branch          32'bxxxxxxxxxxxxxxxxxxxxxxxxx1100011
`define jump            32'bxxxxxxxxxxxxxxxxxxxxxxxxx1100111
`define jalr            32'bxxxxxxxxxxxxxxxxxxxxxxxxx1100111
`define auipc           32'bxxxxxxxxxxxxxxxxxxxxxxxxx0010111
`define lui             32'bxxxxxxxxxxxxxxxxxxxxxxxxx0110111
