`define arithmetic_base 7'b0110011
`define arithmetic_imm  7'b0010011
`define load            7'b0000011
`define store           7'b0100011
`define branch          7'b1100011
`define jump            7'b1101111
`define jalr            7'b1100111
`define auipc           32'bxxxxxxxxxxxxxxxxxxxxxxxxx0010111
`define lui             32'bxxxxxxxxxxxxxxxxxxxxxxxxx0110111
