`define arithmetic      7'b0x10011
`define load            7'b0000011
`define store           7'b0100011
`define branch          7'b1100011
`define jump            7'b1101111
`define jalr            7'b1100111
`define auipc           7'b0010111
`define lui             7'b0110111
