`define ADD 3'b000
`define SUB 3'b001
`define AND 3'b010
`define OR  3'b011
`define XOR 3'b100
`define SLL 3'b101
`define SLR 3'b110
`define SAR 3'b111