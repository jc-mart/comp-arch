// Base ALU ops
`define add 3'b000
`define sub 3'b001
`define and 3'b010
`define or  3'b011
`define xor 3'b100
`define sll 3'b101
`define slr 3'b110
`define sar 3'b111

// ALU input 2 source
`define rf 2'b00
`define se 2'b01
`define ze 2'b10